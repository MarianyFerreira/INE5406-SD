--- Algoritmo para teste do LCD
--- Edson manoel da silva

LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
USE IEEE.NUMERIC_STD.ALL;


ENTITY TESTE_LCD IS
	PORT
		(
		--//	Host Side
		iCLK,iRST_N : IN STD_LOGIC;
		--//	LCD Side
		LCD_DATA : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)	;
		LCD_RW,LCD_EN,LCD_RS : OUT STD_LOGIC
		);
END ENTITY;

ARCHITECTURE FUNCIONAMENTO OF TESTE_LCD IS

SIGNAL LUT_INDEX : STD_LOGIC_VECTOR(5 DOWNTO 0);
SIGNAL LUT_DATA  : STD_LOGIC_VECTOR(8 DOWNTO 0);
SIGNAL mLCD_ST	 : STD_LOGIC_VECTOR(5 DOWNTO 0);
SIGNAL mDLY		 : STD_LOGIC_VECTOR(17 DOWNTO 0);
SIGNAL mLCD_Start: STD_LOGIC;
SIGNAL mLCD_DATA : STD_LOGIC_VECTOR(7 DOWNTO 0);
SIGNAL mLCD_RS	 : STD_LOGIC;
SIGNAL mLCD_Done : STD_LOGIC;

CONSTANT	LCD_INTIAL	: STD_LOGIC_VECTOR(5 DOWNTO 0) := (OTHERS => '0'); --0;
CONSTANT	LCD_LINE1	: STD_LOGIC_VECTOR(5 DOWNTO 0) :=  "000101";	   --5;
CONSTANT	LCD_CH_LINE	: STD_LOGIC_VECTOR(5 DOWNTO 0) :=	LCD_LINE1+ "010000"; --16;
CONSTANT	LCD_LINE2	: STD_LOGIC_VECTOR(5 DOWNTO 0) :=	LCD_LINE1+"010000"+"000001"; --16+1;
CONSTANT	LUT_SIZE	: STD_LOGIC_VECTOR(5 DOWNTO 0) :=	LCD_LINE1+"100000"+"000001";--32+1;


COMPONENT LCD_CONTROLADOR
	PORT
	(
		iDATA		:	 IN STD_LOGIC_VECTOR(7 DOWNTO 0);
		iRS		:	 IN STD_LOGIC;
		iStart		:	 IN STD_LOGIC;
		iCLK		:	 IN STD_LOGIC;
		iRST_N		:	 IN STD_LOGIC;
		oDone		:	 OUT STD_LOGIC;
		LCD_DATA		:	 OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
		LCD_EN		:	 OUT STD_LOGIC;
		LCD_RW		:	 OUT STD_LOGIC;
		LCD_RS		:	 OUT STD_LOGIC
	);
END COMPONENT;


BEGIN


LCDINST:LCD_CONTROLADOR
	PORT MAP
		(	
			--//	Host Side
			iDATA => mLCD_DATA,
			iRS	  => mLCD_RS,
			iStart=> mLCD_Start,
			oDone => mLCD_Done,
			iCLK  => iCLK,
			iRST_N=> iRST_N,
			--//	LCD Interface
			LCD_DATA=>LCD_DATA,
			LCD_RW => LCD_RW,
			LCD_EN => LCD_EN,
			LCD_RS => LCD_RS	
		);

	PROCESS(iCLK,iRST_N)
	BEGIN
		IF(iRST_N = '0') THEN
			LUT_INDEX	<=	(OTHERS => '0');
			mLCD_ST		<=	(OTHERS => '0');
			mDLY		<=	(OTHERS => '0');
			mLCD_Start	<=	'0';
			mLCD_DATA	<=	(OTHERS => '0');
			mLCD_RS		<=	'0';
		ELSIF(iCLK'EVENT AND iCLK = '1') THEN
			IF(LUT_INDEX<LUT_SIZE) THEN
				CASE(mLCD_ST) IS
					WHEN  "000000" =>
						mLCD_DATA	<=	LUT_DATA(7 DOWNTO 0);	-- PASSA O DADO A SER ESCRITO PARA O LCD
						mLCD_RS		<=	LUT_DATA(8);			-- PASSA O SINAL DE RS(DENTRO DO CONTROLADOR ESSE SINAL APENAS É UM BYPASS)
						mLCD_Start	<=	'1';					-- INICIA O LCD
						mLCD_ST		<=	"000001";				-- MUDA DE ESTADO
					WHEN  "000001" =>
						IF(mLCD_Done = '1')	THEN				-- SE O LCD RESPONDE
							mLCD_Start	<=	'0';				-- BAIXA O SINAL DE START
							mLCD_ST		<=	"000010";			-- MUDA O ESTADO			
						END IF;
					WHEN  "000010" =>
						IF(mDLY<"111111111111111110")THEN		-- CONTA ATÉ 262142???
							mDLY	<=	mDLY + '1';
						ELSE
							mDLY	<=	(OTHERS => '0');
							mLCD_ST	<=	"000011";				-- MUDA DE ESTADO
						END IF;
					WHEN  "000011" =>
						LUT_INDEX	<=	LUT_INDEX+'1';			-- MUDA O SÍMBOLO ALFANUMÉRICO A SER ESCRITO?
						mLCD_ST	<=	(OTHERS => '0');
					WHEN OTHERS =>
						mLCD_ST		<=	(OTHERS => '0');
				END CASE;
			END IF;
		END IF;
	END PROCESS;

	PROCESS(LUT_INDEX)
	BEGIN
			CASE(LUT_INDEX) IS -- LUT_DATA É RS & SIMBOLO ASCII. Se RS = 1 Manda escrever um caracter, se igual a 0 é uma instruçao(espaço, limpa, muda o cursor)
			--//	Initial
				WHEN  LCD_INTIAL+"00000" 	   => LUT_DATA	<=	"000111000"; --9'h038; -- 
				WHEN  LCD_INTIAL+"00001" 	   => LUT_DATA	<=	"000001100"; --9'h00C; -- 
				WHEN  LCD_INTIAL+"00010" 	   => LUT_DATA	<=	"000000001"; --9'h001; -- Clear Display(limpa a tela)
				WHEN  LCD_INTIAL+"00011" 	   => LUT_DATA	<=	"000000110"; --9'h006; -- 
				WHEN  LCD_INTIAL+"00100" 	   => LUT_DATA	<=	"010000000"; --9'h080; -- Set DDRAM Adress(seta o endereço da DDRAM do LCD)
--				--//	LINHA 1
				WHEN LCD_LINE1+"00000" =>	LUT_DATA	<=	"100100000"; --9'h120;	-- ESPAÇO EM BRANCO
				WHEN LCD_LINE1+"00001" =>	LUT_DATA	<=	"101001111"; --; Letra O
				WHEN LCD_LINE1+"00010" =>	LUT_DATA	<=	"101111100"; --; Letra L
				WHEN LCD_LINE1+"00011" =>	LUT_DATA	<=	"101100001"; --; LETRA A
				WHEN LCD_LINE1+"00100" =>	LUT_DATA	<=	"100100000"; --9'h120; ESPAÇO EM BRANCO
				WHEN LCD_LINE1+"00101" =>	LUT_DATA	<=	"101001000"; --; LETRA H
				WHEN LCD_LINE1+"00110" =>	LUT_DATA	<=	"101100101"; --; LETRA A
				WHEN LCD_LINE1+"00111" =>	LUT_DATA	<=	"101101110"; --; Letra L
				WHEN LCD_LINE1+"01000" =>	LUT_DATA	<=	"101110010"; --; Letra T
				WHEN LCD_LINE1+"01001" =>	LUT_DATA	<=	"101101001"; --; Letra E
				WHEN LCD_LINE1+"01010" =>	LUT_DATA	<=	"101110001"; --; Letra R
				WHEN LCD_LINE1+"01011" =>	LUT_DATA	<=	"101110101"; --; Letra R
				WHEN LCD_LINE1+"01100" =>	LUT_DATA	<=	"101100101"; --; LETRA A
--				WHEN LCD_LINE1+"00001" =>	LUT_DATA	<=	"101010111"; --9'h157;
--				WHEN LCD_LINE1+"00010" =>	LUT_DATA	<=	"101100101"; --9'h165;
--				WHEN LCD_LINE1+"00011" =>	LUT_DATA	<=	"101101100"; --9'h16C;
--				WHEN LCD_LINE1+"00100" =>	LUT_DATA	<=	"101100011"; --9'h163;
--				WHEN LCD_LINE1+"00101" =>	LUT_DATA	<=	"101101111"; --9'h16F;
--				WHEN LCD_LINE1+"00110" =>	LUT_DATA	<=	"101101101"; --9'h16D;
--				WHEN LCD_LINE1+"00111" =>	LUT_DATA	<=	"101100101"; --9'h165;
--				WHEN LCD_LINE1+"01000" =>	LUT_DATA	<=	"100100000"; --9'h120;
--				WHEN LCD_LINE1+"01001" =>	LUT_DATA	<=	"101110100"; --9'h174;
--				WHEN LCD_LINE1+"01010" =>	LUT_DATA	<=	"101101111"; --9'h16F;
--				WHEN LCD_LINE1+"01011" =>	LUT_DATA	<=	"100100000"; --9'h120;
--				WHEN LCD_LINE1+"01100" =>	LUT_DATA	<=	"101110100"; --9'h174;
--				WHEN LCD_LINE1+"01101" => 	LUT_DATA	<=	"101101000"; --9'h168;
--				WHEN LCD_LINE1+"01110" =>	LUT_DATA	<=	"101100101"; --9'h165;
--				WHEN LCD_LINE1+"01111" =>	LUT_DATA	<=	"100100000"; --9'h120;
--				--//	MUDA DE LINHA
--				WHEN LCD_CH_LINE =>			LUT_DATA	<=	"011000000"; --9'h0C0;
--				--//	LINHA 2
--				WHEN LCD_LINE2+"00000" =>	LUT_DATA	<=	"100100000"; --9'h120;	--
--				WHEN LCD_LINE2+"00001" =>	LUT_DATA	<=	"101000001"; --9'h141;	-- LETRA A
--				WHEN LCD_LINE2+"00010" => 	LUT_DATA	<=	"101101100"; --9'h16C;
--				WHEN LCD_LINE2+"00011" =>	LUT_DATA	<=	"101110100"; --9'h174;
--				WHEN LCD_LINE2+"00100" =>	LUT_DATA	<=	"101100101"; --9'h165;
--				WHEN LCD_LINE2+"00101" =>	LUT_DATA	<=	"101110010"; --9'h172;
--				WHEN LCD_LINE2+"00110" =>	LUT_DATA	<=	"101100001"; --9'h161;
--				WHEN LCD_LINE2+"00111" =>	LUT_DATA	<=	"100100000"; --9'h120;
--				WHEN LCD_LINE2+"01000" =>	LUT_DATA	<=	"101000100"; --9'h144;
--				WHEN LCD_LINE2+"01001" =>	LUT_DATA	<=	"101000101"; --9'h145;
--				WHEN LCD_LINE2+"01010" =>	LUT_DATA	<=	"100110010"; --9'h132;
--				WHEN LCD_LINE2+"01011" =>	LUT_DATA	<=	"110110000"; --9'h1B0;
--				WHEN LCD_LINE2+"01100" =>	LUT_DATA	<=	"100110001"; --9'h131;
--				WHEN LCD_LINE2+"01101" =>	LUT_DATA	<=	"100110001"; --9'h131;
--				WHEN LCD_LINE2+"01110" =>	LUT_DATA	<=	"100110101"; --9'h135;
--				WHEN LCD_LINE2+"01111" =>	LUT_DATA	<=	"100100000"; --9'h120;
				WHEN OTHERS =>				LUT_DATA	<=	"100100000"; --9'h120;
			END CASE;
	END PROCESS;







END ARCHITECTURE;