LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
USE ieee.numeric_std.ALL;

ENTITY RESET_DELAY IS
PORT
	(
		iCLK  : IN STD_LOGIC;
		oRESET: OUT STD_LOGIC
	);
END ENTITY;
		
ARCHITECTURE FUNCIONAMENTO OF RESET_DELAY IS

SIGNAL Cont  : STD_LOGIC_VECTOR(19 DOWNTO 0);


BEGIN

		
		
	PROCESS(iCLK)
	BEGIN
		IF(iCLK'EVENT AND iCLK='1') THEN
			IF(Cont = X"FFFFF")THEN
				oRESET	<=	'1';
			ELSE
				Cont	<=	Cont+1;
				oRESET	<=	'0';
			END IF;
		END IF;
	END PROCESS;
	
END ARCHITECTURE;